module rotateWiring(A, B, clk, rst);
    input clk, rst;
    input [3:0] A [15:0];
    output [3:0] B [15:0];
endmodule

module randomPerm0(A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15);
    input [3:0] A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15;
    output [3:0] B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15;
    assign B_0 = A_10;
    assign B_1 = A_7;
    assign B_2 = A_12;
    assign B_3 = A_6;
    assign B_4 = A_11;
    assign B_5 = A_4;
    assign B_6 = A_13;
    assign B_7 = A_3;
    assign B_8 = A_1;
    assign B_9 = A_15;
    assign B_10 = A_14;
    assign B_11 = A_2;
    assign B_12 = A_9;
    assign B_13 = A_0;
    assign B_14 = A_8;
    assign B_15 = A_5;
endmodule

module randomPerm1(A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15);
    input [3:0] A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15;
    output [3:0] B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15;
    assign B_0 = A_8;
    assign B_1 = A_9;
    assign B_2 = A_3;
    assign B_3 = A_1;
    assign B_4 = A_13;
    assign B_5 = A_12;
    assign B_6 = A_5;
    assign B_7 = A_14;
    assign B_8 = A_2;
    assign B_9 = A_4;
    assign B_10 = A_7;
    assign B_11 = A_6;
    assign B_12 = A_0;
    assign B_13 = A_15;
    assign B_14 = A_11;
    assign B_15 = A_10;
endmodule

module randomPerm2(A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15);
    input [3:0] A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15;
    output [3:0] B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15;
    assign B_0 = A_3;
    assign B_1 = A_0;
    assign B_2 = A_14;
    assign B_3 = A_2;
    assign B_4 = A_1;
    assign B_5 = A_15;
    assign B_6 = A_5;
    assign B_7 = A_6;
    assign B_8 = A_13;
    assign B_9 = A_7;
    assign B_10 = A_11;
    assign B_11 = A_9;
    assign B_12 = A_8;
    assign B_13 = A_4;
    assign B_14 = A_12;
    assign B_15 = A_10;
endmodule

module randomPerm3(A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15);
    input [3:0] A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15;
    output [3:0] B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15;
    assign B_0 = A_7;
    assign B_1 = A_6;
    assign B_2 = A_13;
    assign B_3 = A_4;
    assign B_4 = A_5;
    assign B_5 = A_11;
    assign B_6 = A_8;
    assign B_7 = A_10;
    assign B_8 = A_9;
    assign B_9 = A_1;
    assign B_10 = A_12;
    assign B_11 = A_14;
    assign B_12 = A_15;
    assign B_13 = A_0;
    assign B_14 = A_3;
    assign B_15 = A_2;
endmodule

module randomPerm4(A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15);
    input [3:0] A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15;
    output [3:0] B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15;
    assign B_0 = A_6;
    assign B_1 = A_14;
    assign B_2 = A_12;
    assign B_3 = A_5;
    assign B_4 = A_8;
    assign B_5 = A_9;
    assign B_6 = A_1;
    assign B_7 = A_4;
    assign B_8 = A_10;
    assign B_9 = A_11;
    assign B_10 = A_7;
    assign B_11 = A_0;
    assign B_12 = A_15;
    assign B_13 = A_2;
    assign B_14 = A_13;
    assign B_15 = A_3;
endmodule
module randomPerm5(A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15);
    input [3:0] A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15;
    output [3:0] B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15;
    assign B_0 = A_13;
    assign B_1 = A_3;
    assign B_2 = A_12;
    assign B_3 = A_10;
    assign B_4 = A_5;
    assign B_5 = A_2;
    assign B_6 = A_4;
    assign B_7 = A_7;
    assign B_8 = A_15;
    assign B_9 = A_6;
    assign B_10 = A_1;
    assign B_11 = A_8;
    assign B_12 = A_0;
    assign B_13 = A_9;
    assign B_14 = A_11;
    assign B_15 = A_14;
endmodule
module randomPerm6(A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15);
    input [3:0] A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15;
    output [3:0] B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15;
    assign B_0 = A_12;
    assign B_1 = A_13;
    assign B_2 = A_5;
    assign B_3 = A_0;
    assign B_4 = A_15;
    assign B_5 = A_4;
    assign B_6 = A_1;
    assign B_7 = A_11;
    assign B_8 = A_7;
    assign B_9 = A_6;
    assign B_10 = A_2;
    assign B_11 = A_10;
    assign B_12 = A_14;
    assign B_13 = A_9;
    assign B_14 = A_8;
    assign B_15 = A_3;
endmodule
module randomPerm7(A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15);
    input [3:0] A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15;
    output [3:0] B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7, B_8, B_9, B_10, B_11, B_12, B_13, B_14, B_15;
    assign B_0 = A_5;
    assign B_1 = A_10;
    assign B_2 = A_12;
    assign B_3 = A_11;
    assign B_4 = A_7;
    assign B_5 = A_14;
    assign B_6 = A_6;
    assign B_7 = A_2;
    assign B_8 = A_0;
    assign B_9 = A_4;
    assign B_10 = A_9;
    assign B_11 = A_8;
    assign B_12 = A_15;
    assign B_13 = A_1;
    assign B_14 = A_13;
    assign B_15 = A_3;
endmodule
