module randomPerm3Map(X_all, Y_all, random);
    input [7:0] X_all;
    input random;
    output [7:0] Y_all;
    always @* begin
    
    end
endmodule
